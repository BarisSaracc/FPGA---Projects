----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Baris Sarac
-- 
-- Create Date: 09.09.2025 14:09:21
-- Design Name: 
-- Module Name: COE - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity COE is
--  Port ( );
end COE;

architecture Behavioral of COE is

begin


end Behavioral;
